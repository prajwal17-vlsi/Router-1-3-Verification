package test_pkg;


//import uvm_pkg.sv
	import uvm_pkg::*;
//include uvm_macros.sv
	`include "uvm_macros.svh"
`include "src_xtn.sv"

`include "src_agnt_config.sv"
`include "dst_agnt_config.sv"
`include "env_cfg.sv"

//`include "src_xtn.sv"
`include "src_drv.sv"
`include "src_mon.sv"
`include "src_src_seqr.sv"
`include "src_agnt.sv"
`include "src_agnt_top.sv"
`include "src_src_seqs.sv"

`include "dst_xtn.sv"
//`include "dst_agnt_config.sv"
`include "dst_mon.sv"
`include "dst_seqr.sv"
`include "dst_seqs.sv"
`include "dst_drv.sv"
`include "dst_agnt.sv"
`include "dst_agnt_top.sv"

`include "virtual_sequencer.sv"
`include "virtual_seqs.sv"
`include "sb.sv"

`include "rout_env.sv"


`include "rout_test.sv"
endpackage
